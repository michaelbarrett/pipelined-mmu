MAM�  ��������������٪��������������������������������������˺��˪���������غ�������������������ͩ��������������˹��˩��̺��ݪ��������             Ш      ����    З��    ��ʷ  ����м ����� � ������������а��w�������������	� � ��
�� а   � �     ��A�qb�/��� B��$�Hr#Ǡ$F�Ub$������tu�r1B��>]���<!���<�8.gBh��>;��3��Nx�:��<����:%�:��8�'��_8�v�V;v��{��ޗ����Έ#PΤVо��'�EG���>o.i/B��R�x�5rE�F=}�9�����}/������0��i:@�k.���:�GqFJ@���z8�	�N�W#Ġќ��;��up�|���rF8�8�14�p��ND�PD<����B���0�����|ˮ��p�r���brࣞ�,���8p�k�B'�</��K�����ٮ� �Q9l��{R�y���#��&�(�x��4�_4*E9M����AE���D��2�~so8�ہ�<I������H���|�+��K��Ůx �y.��˰S<X�8�*uH.,�!z$��"���ݣ��Oʋ���6�������Xveϝ�1���V4� $N��8��錛ο7#��S�0�,G��� )0�0��G�`X�g[%��.>�}7j|ԁ5�:�SX���D���(G.X���l���+�g$�?.���X�S~�v�r��d�i�iZ��,�;
��� 
�{�X�a`��~�P�2P���
,l�X��G��;4Y! �`�p����Ĥ�XH��\���(��P`<9�l`P����rk�<���B�.�[��`� SO��|�N*�������_�AοـN��̦~y�1`��'I��vE �~ڦ����[N,٩ (���n�K���� �*�k�cm@b�r�Cu�X�,O��0e �?q �,�5�K��X�Eq��fj�P����tկ��	��2����uS���X�_5���W��A��EɁ�Px~��D0L��i�,tk�U<q"���X��	׀`�������|r=z�P��,��|�?���,20�:Ex��k��X��
,8���w���������%��`u(= ?�l`2�"y@�(׎>0�'�*�0X�N`/�%�����"k�m���u��0�,
[$���N����{�NQ�G^��PC� X#Z�
	$
� �%	*L`d@t|@{������@�CP �#X��G@� �%	*L`d@�|N� b @f~�P6Bp��#XA�HD�@�A%�,��a�2!�	Y>����020?����#���@`A#H�D@�%�,A�	�Lh��0 25z�\�$ڵ���6O�.71�
E�0���$�$A0	JT��&�Fg�|}����D璁�A��@��1`L"�� 	y1O��CG<Gg:j= :�u��j:�����#�H��}�MyzOT��	OoG� ����$9pc�AT�H=`=�9 t����T�$��;n��|.`'O[�P8H?�o1Dn��(��t,^�N�@H��t�{U����X#G�F��D�B�L��gT,�����o=�CT�8��2X��0!��QB����\�G�\�G�\FG
���r:*�:T�Ku��W�Q!W�Q!��Q!�٣B\�G��r�
r���5*���!rQ̭`o���ELE6�4A�`7! A�
���l*$����=T* &j������ʣ��Cs��0��m�<�a�D"(�iF�#������$	&J@X� �о("�%���!��
��1zD@B �%��'"�!U	,|��<R&@�|>p�����������*DB�T�g��#h� 	(It.$VҘ���2��\5CT�\4C��e1T��l�`e �b36@pBQD�B2} �P��QH��F���m {jMp���� bf@�~6PpB��@�"F�8���ghK=�6N�8tN�эN�󋝌�tr�`��(��|Hu@��� ��p���G@`�;�j�����Z2 ���p� :�gx�P��8 �4`|�v�� ہ���<jx�B��,<�/@� ~��!�A[�?(D�$FA#	"I h�OGN ������v��"<,���$�C����M%*�sb����!� DA#	IN{�(�D%�E���΅Ao�6��Y��,��,�(�E`u#E�BѐGBx�nJ�Ә�X���5��@���i�/��@�(�p9�z�t��H^���a0��܀��!0���E�lL��G@� �A%	,L�l�}�0�020P4�U���`�C �@\�"5B!�HD�@�A%	,L�j���?��k�!kA �ą�0CL4?��!
j�!	�X�#	$>�����N?�fsh��5Gp@� �ےih�A��1����c�u1�� p� 0Ġ�e�0x3������w�4�`�c���@9�iق����C�� ��p[�bR!Y	0M�O��[�bXJ � ��l�_� W�"8�*FQ"�ЯS�Wf7B�f��a� [}n���Â�Bp�a�cD�)�"�Xj9b!	�ē$`����	˄W�rm+�`���u0��l���!(��cD1)��Bj�:�pHHDN&a@	�J�&�2VA���Y�1 +Ht�faig��j��nK��t�@��"F�8���
�^D0M�(!P	K`� ��� � P1�n �� �:m���!0��"��JD�#����s�	��	i8G���xL���D�&�!�e�����` b�Zw�f�D4����`�r�tB�(B`�#h� 	�HH�`��%	2>��� �̀�
#D�&82�	A��V�-C�x@:b>�s�aug�C���)u�j�c�;&w0����g8h(��)@8A`���x0=�2A�͹�Fǔ8�:`v���X?+FA{����p���,�fs��jz�|�h:)�����;k����PSA^����v�������^T���������(�� v��r��&��1P�r����y�0 � ����1��L���"|0��hK��`� �CP �#X&K	�Bb�!Un-�	�R���@�&�`	�0���K9#Qx=��������AtA�_|| ~p>�>`>�?�|���A�A��t=(7 _��A���H�W;Ң12H6��؝�UJĮ)�'qSP�	I��� a���5���L4Ҁ}���b��B = i�Q��?z�T�m������	I�@E.#f�r�~0��>*�Z>*�z?*ryh퐃*���1�.i`�i���i��!�#~�vj�!�>�s��3����A�T�gL�<X�2N��A�\0G
�u�T�u����jC.�aw�4�;k�Z�������46�Sna�ׅw;���`A(�,F<��0(SP(Ĕ+t`��Ff��A$H3+0���T��+
t�}�
J�@��6��d}b�4b�0��a-#���B.��
��r�r�r�*�7�L�>�����G��
��E.~���G�
�Ꮕ\�G!��QB.�`[��B�Xȭ}2h��f��cY�	��*�'��8�����`����e\�6$p6�n3��`΁$��g�B4�`J0 5��T�5���o�����)@f��	�D&�� ���80[�C����b�Hf��A����h�	�}px��@�`���B(�/�͂Ԁ���{�r��y8��!S]D��C������ 2P� `��e@p��df�����DЫ�N(W�����h�L#@ 5�����< 3�� ����$��!z�����u�><r�>V�zg���p���y ��OC�� ,cz8o9JCa*��;d:*��v�������8����/���/ �� �8 s��R)$�3Y@{CJ��fܢ��B�8�sY
��梴�n�~���9�z�"���.L��؆� �Z`d �~U@�H�F<�-B��0��`� s��4�"���%�H��@,=�?@h�6(F�{]��4ws�ɹI��y�������P�8��/�%�o�g�_��A����A�A�����=�o���#��Pt�h� v}p�O�����1�}<��pt�}�7��
��N�ׇ:q-��R
�dn�o0$i�J��7�܏"��� �h˛6$Y�
��

��
�V��?�$a���r��\�"[Zt	0�АV �@�e��/A��<���`[�}( 1����A�Yf]����as��͗)&7RKo����BD�BP!��O�6!�A�<��"oH��JL�[��� �k �H��b�G�����=w�@���;�QۻE�!����>@:H�l�P,\1�8t�8�x���;: �L��xz�N1	��@�1�H���7�8�C���u.0@����
?ű��G��fP*p9�o���Fs3�����r�R� C4`ƸX=--4E���ك3����j]�gȡI��p�G@� �@%Z�n�@�B(�`h�#	I P�Bz�)(>�:�| vٹ�o� &�{��$�� ����j�)/A��4���2$��M�&&�4��X�KX�c �G�(6��΁�@�n"a_��#C@�`����c3�A���x, ���p���� ���7!�/ŷ6�B)�o�8 u���!	G �V$
"D�B�A��\�E��v�<��V�1&�쨡��QB/���^�Fz�*�<T�kx�Ћ���V�2���m�6T��Y_nV�-�E&���@�A������r��@&P� :(Y��y�t^Z��!���P���?�h
�BƉ�{H{0m@$D<� %��b�8��+iU� ��AT�`x���;�j������z�SdQ���I+�"a �H����I� ��4T������*I�2l�q���T���.7��@?��!
B/��0Q����

��d `hB@��Q�K#v�+�!�A��1�P٥�`�R�9�B4� �:xOZ8�: w���Xo���B7�!źp�+�m[e�XX8�8P;@w���������,�J�6!`�S�(��!>��.m7�_��A@ ����q�P���y���!C$Ā0�����Q���T����A���X(l��� X���(8�",�-�C��!�	0M��0٭01�4@�6i{ !���&������͖�(�5��xQr�%��A�l���#P�H�R-�����;(}d+�R�?�
| | uP���@�A��^�1a�dAn4��4�v8�8P8L7C����	h}px��@| `�����чcDP������������ �5 �@�g
~S�NJ%�@�H��F����~�-�������T����� cn����<�
���%� �`*��ƈ!8 �4`s����11-��E�~����(7X�,�p�⠣\ q�<\̓�� ��+��W +V�Q�0\H�4Y��	n҄�A���Ԁ�܅�0#V�5��r,�A^�.X0ؤ����c 3�� ��8��n��}ƻ!��hH���P�i��w���������ڽ�pA��آƘ�!�
 	�wA�\j�P�_�aP��`�l�Y͍q�'

��A�Y_P��C<A�
���	����1�Pz�O�b�F����)�j?8ViZ�
�B��,o�� E��l����YA�X���L�Eв#��#��y��%�*�	M��,�@��
�`D(��p�%0v�}� Ld¨���l@��@��"8�xh>�4A��݃�'x���(�]�[�/p�`����HP�r ���A�Ѓ�@v�:X|�i���ꃺ����7E���/*�kਡ��QB/�
�R�
�X�
���zT�u����Q��ףB��B�N�
z��>*��&*���Q���APǆ�xX>x>�?h�<���nл[�b(@f��D�9"P��G<� >������؎��A$	$J0Tn�Dhb���b @���x��%4��Z��l?,���@%i�P �f��KC3�V~6PpB��|`F�4],��C"���HD�@�A&
4��J����Qc�1���jV�;^��kT��QX�A^���#�8�:@uDE��TV�렅a@2='E�L���~O�ӡJ0 5��T�5�_��i�'��0��@�A0 �29�D�:��`:Ah��i@�A���j���/��E��p��@�4pc 3��`΁$��g�D4ҀL�@@5������ L���q Ơ @Af�8g��AL@4��J50� T����5��}@�@/��0h�� @Af�4p� >���h��iP�����w����u�  ���a �� �2��H8(��D��K��a���w��\���/����@(3��`΁$��g�B4�`J0 5��T�5�נ}������ �a�2 ̀6�h�A"�|40� F(�4}���7~ 3�̓����H�s�ū1{ Y�e6���[K���cO��k���4$���sc,��<�`C�]p���A�4�yXe�Rm`n@C�Ǌ<�`�s�P�Kd�����G�iL�d@�|h`� d��\l�0���A�A���� @Ɂ؃��� 䠍�h
�ٰ}�\F��:u���i��P�l���!(��n	E�0�����9LwGqQ���{C��A`�9�s`� ����v�	�oc�#��r
9H�x�	20�yqȺ�C��8t�&v�a����F�d3 vtH�Ra"#Ad�AᒺA�~���	J6!U���	m mV��`�A@(���`�<(t7�@���A���uH��p`��p���҃0��H2#Ȍ&1��h���/Gz8B���4Q\p0Z����r"=n3^d�a'���QeD�1�SQe�� ���Թذ�h���2���`���C�T���d ���V7/Itt�LT%�`5���6��A`��?�A	����Ax�#+Xv?Q7��v���`>4uqXOO�aY}U�dhR>k��hu�78Zxgd9(��U�)ax�b���np�Zd%V��Ō�@y`@��d��EҔ���&aŎ#�})ledJ;2�t�1a`T��e1Oc�!����c痟���A�E�	{��&o�~�X���	nk`�X:��̰N2[�U��b������2�`!�ull���,T;IZ�mŲV�<42����Aaܢ���`�R�n���O��s?.z��$SE�v��|���T1 ?EJ���6�������6�l�*A��!�Tk�O<��)�t���	QP��Ć����ed~c�Ԕ�aֿ�%��J�`J�jo���H U^datP+�ARw��`	���� �$�d� ��P
Id�
�s�1��7޷QU�`���NU:z�	a��� �`���=ֲ��5c�v���%
PB�`���Č����*�M����a:A��`k��D�(bcA7�\�?��mdb
��W~�p^bic��5�s��n*Zd�P�r>~'cZ���:��;@`dB�mY&E�/(/`��
�Y��bY��Xb�۶�$�
`��+�yf���d��Jb���b�.���M�-a���c)汄�n%�%'a�A3��J�[�c̊*S�vd	g�1��(�R'`6;�9!�R��`'�T���/���sŻ����d ��К{�c�%��脵���ݩ*]�b��a�b^��ec��u�9��D��c�`쾬
�!�a��U+7^`u`�� mu��Pe�a��Y�h�_���	�aF! C���?U��S:�`8Z����( A�SU�daS�D#�B�Uld`( �'t1̳���c�R:�b��?�&b�Q��y	1b�n�[�4�l��E�̿�)B/��g�����){;��_����h!�"\p������������$��-�2�Ӽ�恋�.\��ˏ][\��pࢅ:s�����.\x��p����APDw�n?��E.�$fD�g"�0������^����n.\���� ��g��!CU��e2������F�FH�aVC��BT�0��1�U�h�GMFHB!�B�!��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  