entity pmu_testb is
end pmu_testb;

architecture pmu_testb of pmu_testb is
begin

	

end pmu_testb;
