library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;

entity three_stage_pipelined_multimedia_tb is
end three_stage_pipelined_multimedia_tb;