[OPENDOC|Aldec.Hde.HdePlugIn.7|.\pipelined_mmu\src/ib.vhd|]
TemplateId=0
[OPENDOC|Aldec.Hde.HdePlugIn.7|.\pipelined_mmu\src/rf.vhd|]
TemplateId=0
[OPENDOC|Aldec.Hde.HdePlugIn.7|.\pipelined_mmu\src/alu.vhd|]
TemplateId=0
ActiveDocument=1
[OPENDOC|Aldec.Hde.HdePlugIn.7|.\pipelined_mmu\src/decoder.vhd|]
TemplateId=0
[OPENDOC|Aldec.Hde.HdePlugIn.7|.\pipelined_mmu\src/pmu.vhd|]
TemplateId=0
[OPENDOC|Aldec.Hde.HdePlugIn.7|.\pipelined_mmu\src/program_counter.vhd|]
TemplateId=0
[OPENDOC|Aldec.Hde.HdePlugIn.7|.\pipelined_mmu\src/pmu_TB.vhd|]
TemplateId=0
[OPENDOC|Aldec.Hde.HdePlugIn.7|.\pipelined_mmu\src/alu_TB.vhd|]
TemplateId=0
                                                                                                                                                                                                                                                                                                                                                                                                                                                                    