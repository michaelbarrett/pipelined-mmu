[COMPILESTATUS|.\src\ib.vhd]
FileTimeLow=30706295
Status=Modified
[COMPILESTATUS|.\src\rf.vhd]
FileTimeLow=30706295
Status=Modified
[CACHEDOC|Aldec.Project.Generic.7|.\pipelined_mmu\pipelined_mmu.adf|]
Path=
[COMPILESTATUS|.\src\alu.vhd]
FileTimeLow=30706295
Status=Modified
[COMPILESTATUS|.\src\decoder.vhd]
FileTimeLow=30706295
Status=Modified
[COMPILESTATUS|.\src\id_exe_register.vhd]
FileTimeLow=30706142
Status=Compiled
[COMPILESTATUS|.\src\if_id_register.vhd]
FileTimeLow=30706142
Status=Compiled
[COMPILESTATUS|.\src\pmu.vhd]
FileTimeLow=30706295
Status=Modified
[COMPILESTATUS|.\src\pmu_TB.vhd]
FileTimeLow=30706295
Status=Modified
[COMPILESTATUS|.\src\program_counter.vhd]
FileTimeLow=30706295
Status=Modified
[COMPILESTATUS|.\src\alu_TB.vhd]
FileTimeLow=30706295
Status=Modified
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            